//apb slave basic sequence
`include "uvm_macros.svh"
import uvm_pkg::*;

class apb_slave_basic_seq extends uvm_sequence;

endclass
`include "riscv_fetch.sv"
`include "riscv_decode.sv"
`include "riscv_regfile.sv"
`include "riscv_execute.sv"
`include "riscv_dmem.sv"
`include "riscv_control.sv"
module riscv_top(
	input		wire		clk,
	input		wire		reset
);
//TODO: connect and instantiate all sub modules.
endmodule
`include "riscv_fetch.sv"
`include "riscv_decode.sv"

module riscv_top(
	input		wire		clk,
	input		wire		reset
);
//TODO: connect and instantiate all sub modules.
endmodule
//apb slave test
`include "uvm_macros.svh"
import uvm_pkg::*;

class apb_slave_test extends uvm_test;
  
endclass
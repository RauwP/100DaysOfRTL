class day22;

	function new();
	endfunction
	
	function void print_hello();
		$display("Hello, day22 out of #100daysofRTL!");
	endfunction;
endclass
